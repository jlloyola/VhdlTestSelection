library ieee;
  use ieee.std_logic_1164.all;

package PkgAdcFifoConfig is
  constant kAiFifoFullSize : positive := 5;
end PkgAdcFifoConfig;
